
module aes_table3(
                input wire [7 : 0]  tab3_i,
                output wire [31 : 0] tab3_o
               );


  //----------------------------------------------------------------
  // The sbox array.
  //----------------------------------------------------------------
  wire [31 : 0] tab3 [0 : 255];


  //----------------------------------------------------------------
  // Four parallel muxes.
  //----------------------------------------------------------------
  assign tab3_o = tab3[tab3_i];

  assign tab3[8'h00] = 32'h63c6a563;
  assign tab3[8'h01] = 32'h7cf8847c;
  assign tab3[8'h02] = 32'h77ee9977;
  assign tab3[8'h03] = 32'h7bf68d7b;
  assign tab3[8'h04] = 32'hf2ff0df2;
  assign tab3[8'h05] = 32'h6bd6bd6b;
  assign tab3[8'h06] = 32'h6fdeb16f;
  assign tab3[8'h07] = 32'hc59154c5;
  assign tab3[8'h08] = 32'h30605030;
  assign tab3[8'h09] = 32'h01020301;
  assign tab3[8'h0a] = 32'h67cea967;
  assign tab3[8'h0b] = 32'h2b567d2b;
  assign tab3[8'h0c] = 32'hfee719fe;
  assign tab3[8'h0d] = 32'hd7b562d7;
  assign tab3[8'h0e] = 32'hab4de6ab;
  assign tab3[8'h0f] = 32'h76ec9a76;
  assign tab3[8'h10] = 32'hca8f45ca;
  assign tab3[8'h11] = 32'h821f9d82;
  assign tab3[8'h12] = 32'hc98940c9;
  assign tab3[8'h13] = 32'h7dfa877d;
  assign tab3[8'h14] = 32'hfaef15fa;
  assign tab3[8'h15] = 32'h59b2eb59;
  assign tab3[8'h16] = 32'h478ec947;
  assign tab3[8'h17] = 32'hf0fb0bf0;
  assign tab3[8'h18] = 32'had41ecad;
  assign tab3[8'h19] = 32'hd4b367d4;
  assign tab3[8'h1a] = 32'ha25ffda2;
  assign tab3[8'h1b] = 32'haf45eaaf;
  assign tab3[8'h1c] = 32'h9c23bf9c;
  assign tab3[8'h1d] = 32'ha453f7a4;
  assign tab3[8'h1e] = 32'h72e49672;
  assign tab3[8'h1f] = 32'hc09b5bc0;
  assign tab3[8'h20] = 32'hb775c2b7;
  assign tab3[8'h21] = 32'hfde11cfd;
  assign tab3[8'h22] = 32'h933dae93;
  assign tab3[8'h23] = 32'h264c6a26;
  assign tab3[8'h24] = 32'h366c5a36;
  assign tab3[8'h25] = 32'h3f7e413f;
  assign tab3[8'h26] = 32'hf7f502f7;
  assign tab3[8'h27] = 32'hcc834fcc;
  assign tab3[8'h28] = 32'h34685c34;
  assign tab3[8'h29] = 32'ha551f4a5;
  assign tab3[8'h2a] = 32'he5d134e5;
  assign tab3[8'h2b] = 32'hf1f908f1;
  assign tab3[8'h2c] = 32'h71e29371;
  assign tab3[8'h2d] = 32'hd8ab73d8;
  assign tab3[8'h2e] = 32'h31625331;
  assign tab3[8'h2f] = 32'h152a3f15;
  assign tab3[8'h30] = 32'h04080c04;
  assign tab3[8'h31] = 32'hc79552c7;
  assign tab3[8'h32] = 32'h23466523;
  assign tab3[8'h33] = 32'hc39d5ec3;
  assign tab3[8'h34] = 32'h18302818;
  assign tab3[8'h35] = 32'h9637a196;
  assign tab3[8'h36] = 32'h050a0f05;
  assign tab3[8'h37] = 32'h9a2fb59a;
  assign tab3[8'h38] = 32'h070e0907;
  assign tab3[8'h39] = 32'h12243612;
  assign tab3[8'h3a] = 32'h801b9b80;
  assign tab3[8'h3b] = 32'he2df3de2;
  assign tab3[8'h3c] = 32'hebcd26eb;
  assign tab3[8'h3d] = 32'h274e6927;
  assign tab3[8'h3e] = 32'hb27fcdb2;
  assign tab3[8'h3f] = 32'h75ea9f75;
  assign tab3[8'h40] = 32'h09121b09;
  assign tab3[8'h41] = 32'h831d9e83;
  assign tab3[8'h42] = 32'h2c58742c;
  assign tab3[8'h43] = 32'h1a342e1a;
  assign tab3[8'h44] = 32'h1b362d1b;
  assign tab3[8'h45] = 32'h6edcb26e;
  assign tab3[8'h46] = 32'h5ab4ee5a;
  assign tab3[8'h47] = 32'ha05bfba0;
  assign tab3[8'h48] = 32'h52a4f652;
  assign tab3[8'h49] = 32'h3b764d3b;
  assign tab3[8'h4a] = 32'hd6b761d6;
  assign tab3[8'h4b] = 32'hb37dceb3;
  assign tab3[8'h4c] = 32'h29527b29;
  assign tab3[8'h4d] = 32'he3dd3ee3;
  assign tab3[8'h4e] = 32'h2f5e712f;
  assign tab3[8'h4f] = 32'h84139784;
  assign tab3[8'h50] = 32'h53a6f553;
  assign tab3[8'h51] = 32'hd1b968d1;
  assign tab3[8'h52] = 32'h00000000;
  assign tab3[8'h53] = 32'hedc12ced;
  assign tab3[8'h54] = 32'h20406020;
  assign tab3[8'h55] = 32'hfce31ffc;
  assign tab3[8'h56] = 32'hb179c8b1;
  assign tab3[8'h57] = 32'h5bb6ed5b;
  assign tab3[8'h58] = 32'h6ad4be6a;
  assign tab3[8'h59] = 32'hcb8d46cb;
  assign tab3[8'h5a] = 32'hbe67d9be;
  assign tab3[8'h5b] = 32'h39724b39;
  assign tab3[8'h5c] = 32'h4a94de4a;
  assign tab3[8'h5d] = 32'h4c98d44c;
  assign tab3[8'h5e] = 32'h58b0e858;
  assign tab3[8'h5f] = 32'hcf854acf;
  assign tab3[8'h60] = 32'hd0bb6bd0;
  assign tab3[8'h61] = 32'hefc52aef;
  assign tab3[8'h62] = 32'haa4fe5aa;
  assign tab3[8'h63] = 32'hfbed16fb;
  assign tab3[8'h64] = 32'h4386c543;
  assign tab3[8'h65] = 32'h4d9ad74d;
  assign tab3[8'h66] = 32'h33665533;
  assign tab3[8'h67] = 32'h85119485;
  assign tab3[8'h68] = 32'h458acf45;
  assign tab3[8'h69] = 32'hf9e910f9;
  assign tab3[8'h6a] = 32'h02040602;
  assign tab3[8'h6b] = 32'h7ffe817f;
  assign tab3[8'h6c] = 32'h50a0f050;
  assign tab3[8'h6d] = 32'h3c78443c;
  assign tab3[8'h6e] = 32'h9f25ba9f;
  assign tab3[8'h6f] = 32'ha84be3a8;
  assign tab3[8'h70] = 32'h51a2f351;
  assign tab3[8'h71] = 32'ha35dfea3;
  assign tab3[8'h72] = 32'h4080c040;
  assign tab3[8'h73] = 32'h8f058a8f;
  assign tab3[8'h74] = 32'h923fad92;
  assign tab3[8'h75] = 32'h9d21bc9d;
  assign tab3[8'h76] = 32'h38704838;
  assign tab3[8'h77] = 32'hf5f104f5;
  assign tab3[8'h78] = 32'hbc63dfbc;
  assign tab3[8'h79] = 32'hb677c1b6;
  assign tab3[8'h7a] = 32'hdaaf75da;
  assign tab3[8'h7b] = 32'h21426321;
  assign tab3[8'h7c] = 32'h10203010;
  assign tab3[8'h7d] = 32'hffe51aff;
  assign tab3[8'h7e] = 32'hf3fd0ef3;
  assign tab3[8'h7f] = 32'hd2bf6dd2;
  assign tab3[8'h80] = 32'hcd814ccd;
  assign tab3[8'h81] = 32'h0c18140c;
  assign tab3[8'h82] = 32'h13263513;
  assign tab3[8'h83] = 32'hecc32fec;
  assign tab3[8'h84] = 32'h5fbee15f;
  assign tab3[8'h85] = 32'h9735a297;
  assign tab3[8'h86] = 32'h4488cc44;
  assign tab3[8'h87] = 32'h172e3917;
  assign tab3[8'h88] = 32'hc49357c4;
  assign tab3[8'h89] = 32'ha755f2a7;
  assign tab3[8'h8a] = 32'h7efc827e;
  assign tab3[8'h8b] = 32'h3d7a473d;
  assign tab3[8'h8c] = 32'h64c8ac64;
  assign tab3[8'h8d] = 32'h5dbae75d;
  assign tab3[8'h8e] = 32'h19322b19;
  assign tab3[8'h8f] = 32'h73e69573;
  assign tab3[8'h90] = 32'h60c0a060;
  assign tab3[8'h91] = 32'h81199881;
  assign tab3[8'h92] = 32'h4f9ed14f;
  assign tab3[8'h93] = 32'hdca37fdc;
  assign tab3[8'h94] = 32'h22446622;
  assign tab3[8'h95] = 32'h2a547e2a;
  assign tab3[8'h96] = 32'h903bab90;
  assign tab3[8'h97] = 32'h880b8388;
  assign tab3[8'h98] = 32'h468cca46;
  assign tab3[8'h99] = 32'heec729ee;
  assign tab3[8'h9a] = 32'hb86bd3b8;
  assign tab3[8'h9b] = 32'h14283c14;
  assign tab3[8'h9c] = 32'hdea779de;
  assign tab3[8'h9d] = 32'h5ebce25e;
  assign tab3[8'h9e] = 32'h0b161d0b;
  assign tab3[8'h9f] = 32'hdbad76db;
  assign tab3[8'ha0] = 32'he0db3be0;
  assign tab3[8'ha1] = 32'h32645632;
  assign tab3[8'ha2] = 32'h3a744e3a;
  assign tab3[8'ha3] = 32'h0a141e0a;
  assign tab3[8'ha4] = 32'h4992db49;
  assign tab3[8'ha5] = 32'h060c0a06;
  assign tab3[8'ha6] = 32'h24486c24;
  assign tab3[8'ha7] = 32'h5cb8e45c;
  assign tab3[8'ha8] = 32'hc29f5dc2;
  assign tab3[8'ha9] = 32'hd3bd6ed3;
  assign tab3[8'haa] = 32'hac43efac;
  assign tab3[8'hab] = 32'h62c4a662;
  assign tab3[8'hac] = 32'h9139a891;
  assign tab3[8'had] = 32'h9531a495;
  assign tab3[8'hae] = 32'he4d337e4;
  assign tab3[8'haf] = 32'h79f28b79;
  assign tab3[8'hb0] = 32'he7d532e7;
  assign tab3[8'hb1] = 32'hc88b43c8;
  assign tab3[8'hb2] = 32'h376e5937;
  assign tab3[8'hb3] = 32'h6ddab76d;
  assign tab3[8'hb4] = 32'h8d018c8d;
  assign tab3[8'hb5] = 32'hd5b164d5;
  assign tab3[8'hb6] = 32'h4e9cd24e;
  assign tab3[8'hb7] = 32'ha949e0a9;
  assign tab3[8'hb8] = 32'h6cd8b46c;
  assign tab3[8'hb9] = 32'h56acfa56;
  assign tab3[8'hba] = 32'hf4f307f4;
  assign tab3[8'hbb] = 32'heacf25ea;
  assign tab3[8'hbc] = 32'h65caaf65;
  assign tab3[8'hbd] = 32'h7af48e7a;
  assign tab3[8'hbe] = 32'hae47e9ae;
  assign tab3[8'hbf] = 32'h08101808;
  assign tab3[8'hc0] = 32'hba6fd5ba;
  assign tab3[8'hc1] = 32'h78f08878;
  assign tab3[8'hc2] = 32'h254a6f25;
  assign tab3[8'hc3] = 32'h2e5c722e;
  assign tab3[8'hc4] = 32'h1c38241c;
  assign tab3[8'hc5] = 32'ha657f1a6;
  assign tab3[8'hc6] = 32'hb473c7b4;
  assign tab3[8'hc7] = 32'hc69751c6;
  assign tab3[8'hc8] = 32'he8cb23e8;
  assign tab3[8'hc9] = 32'hdda17cdd;
  assign tab3[8'hca] = 32'h74e89c74;
  assign tab3[8'hcb] = 32'h1f3e211f;
  assign tab3[8'hcc] = 32'h4b96dd4b;
  assign tab3[8'hcd] = 32'hbd61dcbd;
  assign tab3[8'hce] = 32'h8b0d868b;
  assign tab3[8'hcf] = 32'h8a0f858a;
  assign tab3[8'hd0] = 32'h70e09070;
  assign tab3[8'hd1] = 32'h3e7c423e;
  assign tab3[8'hd2] = 32'hb571c4b5;
  assign tab3[8'hd3] = 32'h66ccaa66;
  assign tab3[8'hd4] = 32'h4890d848;
  assign tab3[8'hd5] = 32'h03060503;
  assign tab3[8'hd6] = 32'hf6f701f6;
  assign tab3[8'hd7] = 32'h0e1c120e;
  assign tab3[8'hd8] = 32'h61c2a361;
  assign tab3[8'hd9] = 32'h356a5f35;
  assign tab3[8'hda] = 32'h57aef957;
  assign tab3[8'hdb] = 32'hb969d0b9;
  assign tab3[8'hdc] = 32'h86179186;
  assign tab3[8'hdd] = 32'hc19958c1;
  assign tab3[8'hde] = 32'h1d3a271d;
  assign tab3[8'hdf] = 32'h9e27b99e;
  assign tab3[8'he0] = 32'he1d938e1;
  assign tab3[8'he1] = 32'hf8eb13f8;
  assign tab3[8'he2] = 32'h982bb398;
  assign tab3[8'he3] = 32'h11223311;
  assign tab3[8'he4] = 32'h69d2bb69;
  assign tab3[8'he5] = 32'hd9a970d9;
  assign tab3[8'he6] = 32'h8e07898e;
  assign tab3[8'he7] = 32'h9433a794;
  assign tab3[8'he8] = 32'h9b2db69b;
  assign tab3[8'he9] = 32'h1e3c221e;
  assign tab3[8'hea] = 32'h87159287;
  assign tab3[8'heb] = 32'he9c920e9;
  assign tab3[8'hec] = 32'hce8749ce;
  assign tab3[8'hed] = 32'h55aaff55;
  assign tab3[8'hee] = 32'h28507828;
  assign tab3[8'hef] = 32'hdfa57adf;
  assign tab3[8'hf0] = 32'h8c038f8c;
  assign tab3[8'hf1] = 32'ha159f8a1;
  assign tab3[8'hf2] = 32'h89098089;
  assign tab3[8'hf3] = 32'h0d1a170d;
  assign tab3[8'hf4] = 32'hbf65dabf;
  assign tab3[8'hf5] = 32'he6d731e6;
  assign tab3[8'hf6] = 32'h4284c642;
  assign tab3[8'hf7] = 32'h68d0b868;
  assign tab3[8'hf8] = 32'h4182c341;
  assign tab3[8'hf9] = 32'h9929b099;
  assign tab3[8'hfa] = 32'h2d5a772d;
  assign tab3[8'hfb] = 32'h0f1e110f;
  assign tab3[8'hfc] = 32'hb07bcbb0;
  assign tab3[8'hfd] = 32'h54a8fc54;
  assign tab3[8'hfe] = 32'hbb6dd6bb;
  assign tab3[8'hff] = 32'h162c3a16;
  endmodule
