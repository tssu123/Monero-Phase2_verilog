
module aes_table4(
                input wire [7 : 0]  tab4_i,
                output wire [31 : 0] tab4_o
               );


  //----------------------------------------------------------------
  // The sbox array.
  //----------------------------------------------------------------
  wire [31 : 0] tab4 [0 : 255];


  //----------------------------------------------------------------
  // Four parallel muxes.
  //----------------------------------------------------------------
  assign tab4_o = tab4[tab4_i];

  assign tab4[8'h00] = 32'hc6a56363;
  assign tab4[8'h01] = 32'hf8847c7c;
  assign tab4[8'h02] = 32'hee997777;
  assign tab4[8'h03] = 32'hf68d7b7b;
  assign tab4[8'h04] = 32'hff0df2f2;
  assign tab4[8'h05] = 32'hd6bd6b6b;
  assign tab4[8'h06] = 32'hdeb16f6f;
  assign tab4[8'h07] = 32'h9154c5c5;
  assign tab4[8'h08] = 32'h60503030;
  assign tab4[8'h09] = 32'h02030101;
  assign tab4[8'h0a] = 32'hcea96767;
  assign tab4[8'h0b] = 32'h567d2b2b;
  assign tab4[8'h0c] = 32'he719fefe;
  assign tab4[8'h0d] = 32'hb562d7d7;
  assign tab4[8'h0e] = 32'h4de6abab;
  assign tab4[8'h0f] = 32'hec9a7676;
  assign tab4[8'h10] = 32'h8f45caca;
  assign tab4[8'h11] = 32'h1f9d8282;
  assign tab4[8'h12] = 32'h8940c9c9;
  assign tab4[8'h13] = 32'hfa877d7d;
  assign tab4[8'h14] = 32'hef15fafa;
  assign tab4[8'h15] = 32'hb2eb5959;
  assign tab4[8'h16] = 32'h8ec94747;
  assign tab4[8'h17] = 32'hfb0bf0f0;
  assign tab4[8'h18] = 32'h41ecadad;
  assign tab4[8'h19] = 32'hb367d4d4;
  assign tab4[8'h1a] = 32'h5ffda2a2;
  assign tab4[8'h1b] = 32'h45eaafaf;
  assign tab4[8'h1c] = 32'h23bf9c9c;
  assign tab4[8'h1d] = 32'h53f7a4a4;
  assign tab4[8'h1e] = 32'he4967272;
  assign tab4[8'h1f] = 32'h9b5bc0c0;
  assign tab4[8'h20] = 32'h75c2b7b7;
  assign tab4[8'h21] = 32'he11cfdfd;
  assign tab4[8'h22] = 32'h3dae9393;
  assign tab4[8'h23] = 32'h4c6a2626;
  assign tab4[8'h24] = 32'h6c5a3636;
  assign tab4[8'h25] = 32'h7e413f3f;
  assign tab4[8'h26] = 32'hf502f7f7;
  assign tab4[8'h27] = 32'h834fcccc;
  assign tab4[8'h28] = 32'h685c3434;
  assign tab4[8'h29] = 32'h51f4a5a5;
  assign tab4[8'h2a] = 32'hd134e5e5;
  assign tab4[8'h2b] = 32'hf908f1f1;
  assign tab4[8'h2c] = 32'he2937171;
  assign tab4[8'h2d] = 32'hab73d8d8;
  assign tab4[8'h2e] = 32'h62533131;
  assign tab4[8'h2f] = 32'h2a3f1515;
  assign tab4[8'h30] = 32'h080c0404;
  assign tab4[8'h31] = 32'h9552c7c7;
  assign tab4[8'h32] = 32'h46652323;
  assign tab4[8'h33] = 32'h9d5ec3c3;
  assign tab4[8'h34] = 32'h30281818;
  assign tab4[8'h35] = 32'h37a19696;
  assign tab4[8'h36] = 32'h0a0f0505;
  assign tab4[8'h37] = 32'h2fb59a9a;
  assign tab4[8'h38] = 32'h0e090707;
  assign tab4[8'h39] = 32'h24361212;
  assign tab4[8'h3a] = 32'h1b9b8080;
  assign tab4[8'h3b] = 32'hdf3de2e2;
  assign tab4[8'h3c] = 32'hcd26ebeb;
  assign tab4[8'h3d] = 32'h4e692727;
  assign tab4[8'h3e] = 32'h7fcdb2b2;
  assign tab4[8'h3f] = 32'hea9f7575;
  assign tab4[8'h40] = 32'h121b0909;
  assign tab4[8'h41] = 32'h1d9e8383;
  assign tab4[8'h42] = 32'h58742c2c;
  assign tab4[8'h43] = 32'h342e1a1a;
  assign tab4[8'h44] = 32'h362d1b1b;
  assign tab4[8'h45] = 32'hdcb26e6e;
  assign tab4[8'h46] = 32'hb4ee5a5a;
  assign tab4[8'h47] = 32'h5bfba0a0;
  assign tab4[8'h48] = 32'ha4f65252;
  assign tab4[8'h49] = 32'h764d3b3b;
  assign tab4[8'h4a] = 32'hb761d6d6;
  assign tab4[8'h4b] = 32'h7dceb3b3;
  assign tab4[8'h4c] = 32'h527b2929;
  assign tab4[8'h4d] = 32'hdd3ee3e3;
  assign tab4[8'h4e] = 32'h5e712f2f;
  assign tab4[8'h4f] = 32'h13978484;
  assign tab4[8'h50] = 32'ha6f55353;
  assign tab4[8'h51] = 32'hb968d1d1;
  assign tab4[8'h52] = 32'h00000000;
  assign tab4[8'h53] = 32'hc12ceded;
  assign tab4[8'h54] = 32'h40602020;
  assign tab4[8'h55] = 32'he31ffcfc;
  assign tab4[8'h56] = 32'h79c8b1b1;
  assign tab4[8'h57] = 32'hb6ed5b5b;
  assign tab4[8'h58] = 32'hd4be6a6a;
  assign tab4[8'h59] = 32'h8d46cbcb;
  assign tab4[8'h5a] = 32'h67d9bebe;
  assign tab4[8'h5b] = 32'h724b3939;
  assign tab4[8'h5c] = 32'h94de4a4a;
  assign tab4[8'h5d] = 32'h98d44c4c;
  assign tab4[8'h5e] = 32'hb0e85858;
  assign tab4[8'h5f] = 32'h854acfcf;
  assign tab4[8'h60] = 32'hbb6bd0d0;
  assign tab4[8'h61] = 32'hc52aefef;
  assign tab4[8'h62] = 32'h4fe5aaaa;
  assign tab4[8'h63] = 32'hed16fbfb;
  assign tab4[8'h64] = 32'h86c54343;
  assign tab4[8'h65] = 32'h9ad74d4d;
  assign tab4[8'h66] = 32'h66553333;
  assign tab4[8'h67] = 32'h11948585;
  assign tab4[8'h68] = 32'h8acf4545;
  assign tab4[8'h69] = 32'he910f9f9;
  assign tab4[8'h6a] = 32'h04060202;
  assign tab4[8'h6b] = 32'hfe817f7f;
  assign tab4[8'h6c] = 32'ha0f05050;
  assign tab4[8'h6d] = 32'h78443c3c;
  assign tab4[8'h6e] = 32'h25ba9f9f;
  assign tab4[8'h6f] = 32'h4be3a8a8;
  assign tab4[8'h70] = 32'ha2f35151;
  assign tab4[8'h71] = 32'h5dfea3a3;
  assign tab4[8'h72] = 32'h80c04040;
  assign tab4[8'h73] = 32'h058a8f8f;
  assign tab4[8'h74] = 32'h3fad9292;
  assign tab4[8'h75] = 32'h21bc9d9d;
  assign tab4[8'h76] = 32'h70483838;
  assign tab4[8'h77] = 32'hf104f5f5;
  assign tab4[8'h78] = 32'h63dfbcbc;
  assign tab4[8'h79] = 32'h77c1b6b6;
  assign tab4[8'h7a] = 32'haf75dada;
  assign tab4[8'h7b] = 32'h42632121;
  assign tab4[8'h7c] = 32'h20301010;
  assign tab4[8'h7d] = 32'he51affff;
  assign tab4[8'h7e] = 32'hfd0ef3f3;
  assign tab4[8'h7f] = 32'hbf6dd2d2;
  assign tab4[8'h80] = 32'h814ccdcd;
  assign tab4[8'h81] = 32'h18140c0c;
  assign tab4[8'h82] = 32'h26351313;
  assign tab4[8'h83] = 32'hc32fecec;
  assign tab4[8'h84] = 32'hbee15f5f;
  assign tab4[8'h85] = 32'h35a29797;
  assign tab4[8'h86] = 32'h88cc4444;
  assign tab4[8'h87] = 32'h2e391717;
  assign tab4[8'h88] = 32'h9357c4c4;
  assign tab4[8'h89] = 32'h55f2a7a7;
  assign tab4[8'h8a] = 32'hfc827e7e;
  assign tab4[8'h8b] = 32'h7a473d3d;
  assign tab4[8'h8c] = 32'hc8ac6464;
  assign tab4[8'h8d] = 32'hbae75d5d;
  assign tab4[8'h8e] = 32'h322b1919;
  assign tab4[8'h8f] = 32'he6957373;
  assign tab4[8'h90] = 32'hc0a06060;
  assign tab4[8'h91] = 32'h19988181;
  assign tab4[8'h92] = 32'h9ed14f4f;
  assign tab4[8'h93] = 32'ha37fdcdc;
  assign tab4[8'h94] = 32'h44662222;
  assign tab4[8'h95] = 32'h547e2a2a;
  assign tab4[8'h96] = 32'h3bab9090;
  assign tab4[8'h97] = 32'h0b838888;
  assign tab4[8'h98] = 32'h8cca4646;
  assign tab4[8'h99] = 32'hc729eeee;
  assign tab4[8'h9a] = 32'h6bd3b8b8;
  assign tab4[8'h9b] = 32'h283c1414;
  assign tab4[8'h9c] = 32'ha779dede;
  assign tab4[8'h9d] = 32'hbce25e5e;
  assign tab4[8'h9e] = 32'h161d0b0b;
  assign tab4[8'h9f] = 32'had76dbdb;
  assign tab4[8'ha0] = 32'hdb3be0e0;
  assign tab4[8'ha1] = 32'h64563232;
  assign tab4[8'ha2] = 32'h744e3a3a;
  assign tab4[8'ha3] = 32'h141e0a0a;
  assign tab4[8'ha4] = 32'h92db4949;
  assign tab4[8'ha5] = 32'h0c0a0606;
  assign tab4[8'ha6] = 32'h486c2424;
  assign tab4[8'ha7] = 32'hb8e45c5c;
  assign tab4[8'ha8] = 32'h9f5dc2c2;
  assign tab4[8'ha9] = 32'hbd6ed3d3;
  assign tab4[8'haa] = 32'h43efacac;
  assign tab4[8'hab] = 32'hc4a66262;
  assign tab4[8'hac] = 32'h39a89191;
  assign tab4[8'had] = 32'h31a49595;
  assign tab4[8'hae] = 32'hd337e4e4;
  assign tab4[8'haf] = 32'hf28b7979;
  assign tab4[8'hb0] = 32'hd532e7e7;
  assign tab4[8'hb1] = 32'h8b43c8c8;
  assign tab4[8'hb2] = 32'h6e593737;
  assign tab4[8'hb3] = 32'hdab76d6d;
  assign tab4[8'hb4] = 32'h018c8d8d;
  assign tab4[8'hb5] = 32'hb164d5d5;
  assign tab4[8'hb6] = 32'h9cd24e4e;
  assign tab4[8'hb7] = 32'h49e0a9a9;
  assign tab4[8'hb8] = 32'hd8b46c6c;
  assign tab4[8'hb9] = 32'hacfa5656;
  assign tab4[8'hba] = 32'hf307f4f4;
  assign tab4[8'hbb] = 32'hcf25eaea;
  assign tab4[8'hbc] = 32'hcaaf6565;
  assign tab4[8'hbd] = 32'hf48e7a7a;
  assign tab4[8'hbe] = 32'h47e9aeae;
  assign tab4[8'hbf] = 32'h10180808;
  assign tab4[8'hc0] = 32'h6fd5baba;
  assign tab4[8'hc1] = 32'hf0887878;
  assign tab4[8'hc2] = 32'h4a6f2525;
  assign tab4[8'hc3] = 32'h5c722e2e;
  assign tab4[8'hc4] = 32'h38241c1c;
  assign tab4[8'hc5] = 32'h57f1a6a6;
  assign tab4[8'hc6] = 32'h73c7b4b4;
  assign tab4[8'hc7] = 32'h9751c6c6;
  assign tab4[8'hc8] = 32'hcb23e8e8;
  assign tab4[8'hc9] = 32'ha17cdddd;
  assign tab4[8'hca] = 32'he89c7474;
  assign tab4[8'hcb] = 32'h3e211f1f;
  assign tab4[8'hcc] = 32'h96dd4b4b;
  assign tab4[8'hcd] = 32'h61dcbdbd;
  assign tab4[8'hce] = 32'h0d868b8b;
  assign tab4[8'hcf] = 32'h0f858a8a;
  assign tab4[8'hd0] = 32'he0907070;
  assign tab4[8'hd1] = 32'h7c423e3e;
  assign tab4[8'hd2] = 32'h71c4b5b5;
  assign tab4[8'hd3] = 32'hccaa6666;
  assign tab4[8'hd4] = 32'h90d84848;
  assign tab4[8'hd5] = 32'h06050303;
  assign tab4[8'hd6] = 32'hf701f6f6;
  assign tab4[8'hd7] = 32'h1c120e0e;
  assign tab4[8'hd8] = 32'hc2a36161;
  assign tab4[8'hd9] = 32'h6a5f3535;
  assign tab4[8'hda] = 32'haef95757;
  assign tab4[8'hdb] = 32'h69d0b9b9;
  assign tab4[8'hdc] = 32'h17918686;
  assign tab4[8'hdd] = 32'h9958c1c1;
  assign tab4[8'hde] = 32'h3a271d1d;
  assign tab4[8'hdf] = 32'h27b99e9e;
  assign tab4[8'he0] = 32'hd938e1e1;
  assign tab4[8'he1] = 32'heb13f8f8;
  assign tab4[8'he2] = 32'h2bb39898;
  assign tab4[8'he3] = 32'h22331111;
  assign tab4[8'he4] = 32'hd2bb6969;
  assign tab4[8'he5] = 32'ha970d9d9;
  assign tab4[8'he6] = 32'h07898e8e;
  assign tab4[8'he7] = 32'h33a79494;
  assign tab4[8'he8] = 32'h2db69b9b;
  assign tab4[8'he9] = 32'h3c221e1e;
  assign tab4[8'hea] = 32'h15928787;
  assign tab4[8'heb] = 32'hc920e9e9;
  assign tab4[8'hec] = 32'h8749cece;
  assign tab4[8'hed] = 32'haaff5555;
  assign tab4[8'hee] = 32'h50782828;
  assign tab4[8'hef] = 32'ha57adfdf;
  assign tab4[8'hf0] = 32'h038f8c8c;
  assign tab4[8'hf1] = 32'h59f8a1a1;
  assign tab4[8'hf2] = 32'h09808989;
  assign tab4[8'hf3] = 32'h1a170d0d;
  assign tab4[8'hf4] = 32'h65dabfbf;
  assign tab4[8'hf5] = 32'hd731e6e6;
  assign tab4[8'hf6] = 32'h84c64242;
  assign tab4[8'hf7] = 32'hd0b86868;
  assign tab4[8'hf8] = 32'h82c34141;
  assign tab4[8'hf9] = 32'h29b09999;
  assign tab4[8'hfa] = 32'h5a772d2d;
  assign tab4[8'hfb] = 32'h1e110f0f;
  assign tab4[8'hfc] = 32'h7bcbb0b0;
  assign tab4[8'hfd] = 32'ha8fc5454;
  assign tab4[8'hfe] = 32'h6dd6bbbb;
  assign tab4[8'hff] = 32'h2c3a1616;
  endmodule

