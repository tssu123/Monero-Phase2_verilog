
module aes_table2(
                input wire [7 : 0]  tab2_i,
                output wire [31 : 0] tab2_o
               );


  //----------------------------------------------------------------
  // The sbox array.
  //----------------------------------------------------------------
  wire [31 : 0] tab2 [0 : 255];


  //----------------------------------------------------------------
  // Four parallel muxes.
  //----------------------------------------------------------------
  assign tab2_o = tab2[tab2_i];

  assign tab2[8'h00] = 32'h6363c6a5;
  assign tab2[8'h01] = 32'h7c7cf884;
  assign tab2[8'h02] = 32'h7777ee99;
  assign tab2[8'h03] = 32'h7b7bf68d;
  assign tab2[8'h04] = 32'hf2f2ff0d;
  assign tab2[8'h05] = 32'h6b6bd6bd;
  assign tab2[8'h06] = 32'h6f6fdeb1;
  assign tab2[8'h07] = 32'hc5c59154;
  assign tab2[8'h08] = 32'h30306050;
  assign tab2[8'h09] = 32'h01010203;
  assign tab2[8'h0a] = 32'h6767cea9;
  assign tab2[8'h0b] = 32'h2b2b567d;
  assign tab2[8'h0c] = 32'hfefee719;
  assign tab2[8'h0d] = 32'hd7d7b562;
  assign tab2[8'h0e] = 32'habab4de6;
  assign tab2[8'h0f] = 32'h7676ec9a;
  assign tab2[8'h10] = 32'hcaca8f45;
  assign tab2[8'h11] = 32'h82821f9d;
  assign tab2[8'h12] = 32'hc9c98940;
  assign tab2[8'h13] = 32'h7d7dfa87;
  assign tab2[8'h14] = 32'hfafaef15;
  assign tab2[8'h15] = 32'h5959b2eb;
  assign tab2[8'h16] = 32'h47478ec9;
  assign tab2[8'h17] = 32'hf0f0fb0b;
  assign tab2[8'h18] = 32'hadad41ec;
  assign tab2[8'h19] = 32'hd4d4b367;
  assign tab2[8'h1a] = 32'ha2a25ffd;
  assign tab2[8'h1b] = 32'hafaf45ea;
  assign tab2[8'h1c] = 32'h9c9c23bf;
  assign tab2[8'h1d] = 32'ha4a453f7;
  assign tab2[8'h1e] = 32'h7272e496;
  assign tab2[8'h1f] = 32'hc0c09b5b;
  assign tab2[8'h20] = 32'hb7b775c2;
  assign tab2[8'h21] = 32'hfdfde11c;
  assign tab2[8'h22] = 32'h93933dae;
  assign tab2[8'h23] = 32'h26264c6a;
  assign tab2[8'h24] = 32'h36366c5a;
  assign tab2[8'h25] = 32'h3f3f7e41;
  assign tab2[8'h26] = 32'hf7f7f502;
  assign tab2[8'h27] = 32'hcccc834f;
  assign tab2[8'h28] = 32'h3434685c;
  assign tab2[8'h29] = 32'ha5a551f4;
  assign tab2[8'h2a] = 32'he5e5d134;
  assign tab2[8'h2b] = 32'hf1f1f908;
  assign tab2[8'h2c] = 32'h7171e293;
  assign tab2[8'h2d] = 32'hd8d8ab73;
  assign tab2[8'h2e] = 32'h31316253;
  assign tab2[8'h2f] = 32'h15152a3f;
  assign tab2[8'h30] = 32'h0404080c;
  assign tab2[8'h31] = 32'hc7c79552;
  assign tab2[8'h32] = 32'h23234665;
  assign tab2[8'h33] = 32'hc3c39d5e;
  assign tab2[8'h34] = 32'h18183028;
  assign tab2[8'h35] = 32'h969637a1;
  assign tab2[8'h36] = 32'h05050a0f;
  assign tab2[8'h37] = 32'h9a9a2fb5;
  assign tab2[8'h38] = 32'h07070e09;
  assign tab2[8'h39] = 32'h12122436;
  assign tab2[8'h3a] = 32'h80801b9b;
  assign tab2[8'h3b] = 32'he2e2df3d;
  assign tab2[8'h3c] = 32'hebebcd26;
  assign tab2[8'h3d] = 32'h27274e69;
  assign tab2[8'h3e] = 32'hb2b27fcd;
  assign tab2[8'h3f] = 32'h7575ea9f;
  assign tab2[8'h40] = 32'h0909121b;
  assign tab2[8'h41] = 32'h83831d9e;
  assign tab2[8'h42] = 32'h2c2c5874;
  assign tab2[8'h43] = 32'h1a1a342e;
  assign tab2[8'h44] = 32'h1b1b362d;
  assign tab2[8'h45] = 32'h6e6edcb2;
  assign tab2[8'h46] = 32'h5a5ab4ee;
  assign tab2[8'h47] = 32'ha0a05bfb;
  assign tab2[8'h48] = 32'h5252a4f6;
  assign tab2[8'h49] = 32'h3b3b764d;
  assign tab2[8'h4a] = 32'hd6d6b761;
  assign tab2[8'h4b] = 32'hb3b37dce;
  assign tab2[8'h4c] = 32'h2929527b;
  assign tab2[8'h4d] = 32'he3e3dd3e;
  assign tab2[8'h4e] = 32'h2f2f5e71;
  assign tab2[8'h4f] = 32'h84841397;
  assign tab2[8'h50] = 32'h5353a6f5;
  assign tab2[8'h51] = 32'hd1d1b968;
  assign tab2[8'h52] = 32'h00000000;
  assign tab2[8'h53] = 32'hededc12c;
  assign tab2[8'h54] = 32'h20204060;
  assign tab2[8'h55] = 32'hfcfce31f;
  assign tab2[8'h56] = 32'hb1b179c8;
  assign tab2[8'h57] = 32'h5b5bb6ed;
  assign tab2[8'h58] = 32'h6a6ad4be;
  assign tab2[8'h59] = 32'hcbcb8d46;
  assign tab2[8'h5a] = 32'hbebe67d9;
  assign tab2[8'h5b] = 32'h3939724b;
  assign tab2[8'h5c] = 32'h4a4a94de;
  assign tab2[8'h5d] = 32'h4c4c98d4;
  assign tab2[8'h5e] = 32'h5858b0e8;
  assign tab2[8'h5f] = 32'hcfcf854a;
  assign tab2[8'h60] = 32'hd0d0bb6b;
  assign tab2[8'h61] = 32'hefefc52a;
  assign tab2[8'h62] = 32'haaaa4fe5;
  assign tab2[8'h63] = 32'hfbfbed16;
  assign tab2[8'h64] = 32'h434386c5;
  assign tab2[8'h65] = 32'h4d4d9ad7;
  assign tab2[8'h66] = 32'h33336655;
  assign tab2[8'h67] = 32'h85851194;
  assign tab2[8'h68] = 32'h45458acf;
  assign tab2[8'h69] = 32'hf9f9e910;
  assign tab2[8'h6a] = 32'h02020406;
  assign tab2[8'h6b] = 32'h7f7ffe81;
  assign tab2[8'h6c] = 32'h5050a0f0;
  assign tab2[8'h6d] = 32'h3c3c7844;
  assign tab2[8'h6e] = 32'h9f9f25ba;
  assign tab2[8'h6f] = 32'ha8a84be3;
  assign tab2[8'h70] = 32'h5151a2f3;
  assign tab2[8'h71] = 32'ha3a35dfe;
  assign tab2[8'h72] = 32'h404080c0;
  assign tab2[8'h73] = 32'h8f8f058a;
  assign tab2[8'h74] = 32'h92923fad;
  assign tab2[8'h75] = 32'h9d9d21bc;
  assign tab2[8'h76] = 32'h38387048;
  assign tab2[8'h77] = 32'hf5f5f104;
  assign tab2[8'h78] = 32'hbcbc63df;
  assign tab2[8'h79] = 32'hb6b677c1;
  assign tab2[8'h7a] = 32'hdadaaf75;
  assign tab2[8'h7b] = 32'h21214263;
  assign tab2[8'h7c] = 32'h10102030;
  assign tab2[8'h7d] = 32'hffffe51a;
  assign tab2[8'h7e] = 32'hf3f3fd0e;
  assign tab2[8'h7f] = 32'hd2d2bf6d;
  assign tab2[8'h80] = 32'hcdcd814c;
  assign tab2[8'h81] = 32'h0c0c1814;
  assign tab2[8'h82] = 32'h13132635;
  assign tab2[8'h83] = 32'hececc32f;
  assign tab2[8'h84] = 32'h5f5fbee1;
  assign tab2[8'h85] = 32'h979735a2;
  assign tab2[8'h86] = 32'h444488cc;
  assign tab2[8'h87] = 32'h17172e39;
  assign tab2[8'h88] = 32'hc4c49357;
  assign tab2[8'h89] = 32'ha7a755f2;
  assign tab2[8'h8a] = 32'h7e7efc82;
  assign tab2[8'h8b] = 32'h3d3d7a47;
  assign tab2[8'h8c] = 32'h6464c8ac;
  assign tab2[8'h8d] = 32'h5d5dbae7;
  assign tab2[8'h8e] = 32'h1919322b;
  assign tab2[8'h8f] = 32'h7373e695;
  assign tab2[8'h90] = 32'h6060c0a0;
  assign tab2[8'h91] = 32'h81811998;
  assign tab2[8'h92] = 32'h4f4f9ed1;
  assign tab2[8'h93] = 32'hdcdca37f;
  assign tab2[8'h94] = 32'h22224466;
  assign tab2[8'h95] = 32'h2a2a547e;
  assign tab2[8'h96] = 32'h90903bab;
  assign tab2[8'h97] = 32'h88880b83;
  assign tab2[8'h98] = 32'h46468cca;
  assign tab2[8'h99] = 32'heeeec729;
  assign tab2[8'h9a] = 32'hb8b86bd3;
  assign tab2[8'h9b] = 32'h1414283c;
  assign tab2[8'h9c] = 32'hdedea779;
  assign tab2[8'h9d] = 32'h5e5ebce2;
  assign tab2[8'h9e] = 32'h0b0b161d;
  assign tab2[8'h9f] = 32'hdbdbad76;
  assign tab2[8'ha0] = 32'he0e0db3b;
  assign tab2[8'ha1] = 32'h32326456;
  assign tab2[8'ha2] = 32'h3a3a744e;
  assign tab2[8'ha3] = 32'h0a0a141e;
  assign tab2[8'ha4] = 32'h494992db;
  assign tab2[8'ha5] = 32'h06060c0a;
  assign tab2[8'ha6] = 32'h2424486c;
  assign tab2[8'ha7] = 32'h5c5cb8e4;
  assign tab2[8'ha8] = 32'hc2c29f5d;
  assign tab2[8'ha9] = 32'hd3d3bd6e;
  assign tab2[8'haa] = 32'hacac43ef;
  assign tab2[8'hab] = 32'h6262c4a6;
  assign tab2[8'hac] = 32'h919139a8;
  assign tab2[8'had] = 32'h959531a4;
  assign tab2[8'hae] = 32'he4e4d337;
  assign tab2[8'haf] = 32'h7979f28b;
  assign tab2[8'hb0] = 32'he7e7d532;
  assign tab2[8'hb1] = 32'hc8c88b43;
  assign tab2[8'hb2] = 32'h37376e59;
  assign tab2[8'hb3] = 32'h6d6ddab7;
  assign tab2[8'hb4] = 32'h8d8d018c;
  assign tab2[8'hb5] = 32'hd5d5b164;
  assign tab2[8'hb6] = 32'h4e4e9cd2;
  assign tab2[8'hb7] = 32'ha9a949e0;
  assign tab2[8'hb8] = 32'h6c6cd8b4;
  assign tab2[8'hb9] = 32'h5656acfa;
  assign tab2[8'hba] = 32'hf4f4f307;
  assign tab2[8'hbb] = 32'heaeacf25;
  assign tab2[8'hbc] = 32'h6565caaf;
  assign tab2[8'hbd] = 32'h7a7af48e;
  assign tab2[8'hbe] = 32'haeae47e9;
  assign tab2[8'hbf] = 32'h08081018;
  assign tab2[8'hc0] = 32'hbaba6fd5;
  assign tab2[8'hc1] = 32'h7878f088;
  assign tab2[8'hc2] = 32'h25254a6f;
  assign tab2[8'hc3] = 32'h2e2e5c72;
  assign tab2[8'hc4] = 32'h1c1c3824;
  assign tab2[8'hc5] = 32'ha6a657f1;
  assign tab2[8'hc6] = 32'hb4b473c7;
  assign tab2[8'hc7] = 32'hc6c69751;
  assign tab2[8'hc8] = 32'he8e8cb23;
  assign tab2[8'hc9] = 32'hdddda17c;
  assign tab2[8'hca] = 32'h7474e89c;
  assign tab2[8'hcb] = 32'h1f1f3e21;
  assign tab2[8'hcc] = 32'h4b4b96dd;
  assign tab2[8'hcd] = 32'hbdbd61dc;
  assign tab2[8'hce] = 32'h8b8b0d86;
  assign tab2[8'hcf] = 32'h8a8a0f85;
  assign tab2[8'hd0] = 32'h7070e090;
  assign tab2[8'hd1] = 32'h3e3e7c42;
  assign tab2[8'hd2] = 32'hb5b571c4;
  assign tab2[8'hd3] = 32'h6666ccaa;
  assign tab2[8'hd4] = 32'h484890d8;
  assign tab2[8'hd5] = 32'h03030605;
  assign tab2[8'hd6] = 32'hf6f6f701;
  assign tab2[8'hd7] = 32'h0e0e1c12;
  assign tab2[8'hd8] = 32'h6161c2a3;
  assign tab2[8'hd9] = 32'h35356a5f;
  assign tab2[8'hda] = 32'h5757aef9;
  assign tab2[8'hdb] = 32'hb9b969d0;
  assign tab2[8'hdc] = 32'h86861791;
  assign tab2[8'hdd] = 32'hc1c19958;
  assign tab2[8'hde] = 32'h1d1d3a27;
  assign tab2[8'hdf] = 32'h9e9e27b9;
  assign tab2[8'he0] = 32'he1e1d938;
  assign tab2[8'he1] = 32'hf8f8eb13;
  assign tab2[8'he2] = 32'h98982bb3;
  assign tab2[8'he3] = 32'h11112233;
  assign tab2[8'he4] = 32'h6969d2bb;
  assign tab2[8'he5] = 32'hd9d9a970;
  assign tab2[8'he6] = 32'h8e8e0789;
  assign tab2[8'he7] = 32'h949433a7;
  assign tab2[8'he8] = 32'h9b9b2db6;
  assign tab2[8'he9] = 32'h1e1e3c22;
  assign tab2[8'hea] = 32'h87871592;
  assign tab2[8'heb] = 32'he9e9c920;
  assign tab2[8'hec] = 32'hcece8749;
  assign tab2[8'hed] = 32'h5555aaff;
  assign tab2[8'hee] = 32'h28285078;
  assign tab2[8'hef] = 32'hdfdfa57a;
  assign tab2[8'hf0] = 32'h8c8c038f;
  assign tab2[8'hf1] = 32'ha1a159f8;
  assign tab2[8'hf2] = 32'h89890980;
  assign tab2[8'hf3] = 32'h0d0d1a17;
  assign tab2[8'hf4] = 32'hbfbf65da;
  assign tab2[8'hf5] = 32'he6e6d731;
  assign tab2[8'hf6] = 32'h424284c6;
  assign tab2[8'hf7] = 32'h6868d0b8;
  assign tab2[8'hf8] = 32'h414182c3;
  assign tab2[8'hf9] = 32'h999929b0;
  assign tab2[8'hfa] = 32'h2d2d5a77;
  assign tab2[8'hfb] = 32'h0f0f1e11;
  assign tab2[8'hfc] = 32'hb0b07bcb;
  assign tab2[8'hfd] = 32'h5454a8fc;
  assign tab2[8'hfe] = 32'hbbbb6dd6;
  assign tab2[8'hff] = 32'h16162c3a;
  endmodule	
